    Mac OS X            	   2  �     �                                    ATTR;���  �   �   �                  �   :  com.apple.quarantine   *   �  "com.apple.LaunchServices.OpenWith -7B  �     com.apple.lastuseddate#PS D310081;5c5301cd;Firefox;BC1C779E-E8D7-4D31-987C-7B35E24AE4E0bplist00�WversionTpath_bundleidentifier _$/Applications/Visual Studio Code.app_com.microsoft.VSCode/1X                            o��\    ;T                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    This resource fork intentionally left blank                                                                                                                                                                                                                            ��